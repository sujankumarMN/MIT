//package file
package my_package;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "mul_test.svh"		
endpackage:my_package

