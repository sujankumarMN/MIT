module what(intf i);
endmodule
