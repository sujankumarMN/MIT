package my_pkg;
	`include "uvm_macros.svh"
	import uvm_pkg::*;
	`include "environment.svh"
	`include "test.svh"
endpackage:my_pkg
