class A;
	function new();
		$display("this is 
