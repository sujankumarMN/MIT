
package pack;
`include "uvm_macros.svh"
import uvm_pkg::*;
`include "test.svh"
endpackage

