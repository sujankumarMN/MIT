interface uvm_interface();

endinterface
